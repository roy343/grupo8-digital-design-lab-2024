module BattleshipMain(

	input logic clk,
	output logic hSync,vSync,syncBlank,bSync,
	output logic [7:0]red,green,blue,
	output logic clk25

);

	logic [49:0][9:0] matrix = '{
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
	 {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011},
    {4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0000, 4'b0001, 4'b0010, 4'b0011,4'b0011}
};



	VGAMain VGA(
	clk,
	matrix,
	hSync,
	vSync,
	syncBlank,
	bSync,
	red,
	green,
	blue,
	clk25);
	
endmodule