library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
entity Sumador4bits is
 Port ( A : in STD_LOGIC;
 B : in STD_LOGIC;
 CarryIn : in STD_LOGIC;
 Sum : out STD_LOGIC;
 CarryOut : out STD_LOGIC);
end Sumador4bits;
 
architecture gate of Sumador4bits is
 
begin
 
 
end gate;