
					  