module CheckPos( input logic [9:0] sincronización_horizontal,sincronización_vertical,
					  output logic [24:0]pos);
					  

					  
					  
endmodule
					  