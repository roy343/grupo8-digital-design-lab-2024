module ALU (
    input logic [31:0] A,
    input logic [31:0] B,
    input logic [3:0] opcode,
    output logic [31:0] result,
	 output logic [3:0] ALUFlags
);

    logic [32:0] temp_result; 
	 
	 logic N, Z, C, V 

    always_comb begin
        result = 0;
        N = 0;
        Z = 0;
        C = 0;
        V = 0;

        case(opcode)
            4'b0000: begin // AND
                result = A & B;
            end
            4'b0001: begin // OR
                result = A | B;
            end
            4'b0010: begin // ADD
                temp_result = A + B;
                result = temp_result[31:0];
                C = temp_result[32]; 
                V = (A[31] == B[31]) && (result[31] != A[31]); 
            end
            4'b0011: begin // Multiplication
                result = A * B;
            end
            4'b0100: begin // Division
                result = A / B;
            end
            4'b0101: begin // Modulo
                result = A % B;
            end
            4'b0110: begin // SUB
                temp_result = A - B;
                result = temp_result[31:0];
                C = temp_result[32]; 
                V = (A[31] != B[31]) && (result[31] != A[31]); 
            end
            4'b0111: begin // Shift left
                result = A << B;
            end
            4'b1000: begin // Shift right
                result = A >> B;
            end
            4'b1001: begin // XOR
                result = A ^ B;
            end
            default: begin
                result = 0;
            end
        endcase

        
        N = result[31]; 
        Z = (result == 0); 
    end
	 
	 assign ALUFlags = {N, Z, C, V}
endmodule